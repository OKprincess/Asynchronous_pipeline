// ===================================================
//	=================[ VLSISYS Lab. ]=================
//	* Author		: oksj (oksj@sookmyung.ac.kr)
//	* Filename		: click_network.v
//	* Description	: 
// ===================================================
`include	"click_reg.v"
`include	"click_sink.v"
`include	"click_source.v"

module click_network 
(
	output
);
	
endmodule
